----------------------------------------------------------------------------------
--  This file is part of the ASTERICS Framework.
--  ASTERICS is (C) Hochschule Augsburg, University of Applied Sciences.
----------------------------------------------------------------------------------
-- File:           AXI_Master.vhd
-- Entity:         AXI_Master
--
-- Company:        University of Applied Sciences, Augsburg, Germany
-- Author:         Alexander Zoellner, Michael Schaeferling
--
-- Version:  1.0
-- Modified:
--
-- Description:    An AXI-Master implementation.
-- Comment:        This files content was generated by the Xilinx 
--                 IP Wizard and modified to build an encapsulated 
--                 AXI-Master interface.
----------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;


library axi_master_burst_v2_0_7;
use axi_master_burst_v2_0_7.axi_master_burst;


entity AXI_Master is
  generic
  (
    C_FAMILY                       : string               := "zynq";
    C_M_AXI_ADDR_WIDTH             : integer              := 32;
    C_M_AXI_DATA_WIDTH             : integer              := 32;
    C_MAX_BURST_LEN                : integer              := 16;
    C_NATIVE_DATA_WIDTH            : integer              := 32;
    C_LENGTH_WIDTH                 : integer              := 12;
    C_ADDR_PIPE_DEPTH              : integer              := 1
  );
  port
  (
    -- AXI Master Bus Signals:
    m_axi_aclk                     : in  std_logic;
    m_axi_aresetn                  : in  std_logic;
    md_error                       : out std_logic;
    m_axi_arready                  : in  std_logic;
    m_axi_arvalid                  : out std_logic;
    m_axi_araddr                   : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
    m_axi_arlen                    : out std_logic_vector(7 downto 0);
    m_axi_arsize                   : out std_logic_vector(2 downto 0);
    m_axi_arburst                  : out std_logic_vector(1 downto 0);
    m_axi_arprot                   : out std_logic_vector(2 downto 0);
    m_axi_arcache                  : out std_logic_vector(3 downto 0);
    m_axi_rready                   : out std_logic;
    m_axi_rvalid                   : in  std_logic;
    m_axi_rdata                    : in  std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
    m_axi_rresp                    : in  std_logic_vector(1 downto 0);
    m_axi_rlast                    : in  std_logic;
    m_axi_awready                  : in  std_logic;
    m_axi_awvalid                  : out std_logic;
    m_axi_awaddr                   : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
    m_axi_awlen                    : out std_logic_vector(7 downto 0);
    m_axi_awsize                   : out std_logic_vector(2 downto 0);
    m_axi_awburst                  : out std_logic_vector(1 downto 0);
    m_axi_awprot                   : out std_logic_vector(2 downto 0);
    m_axi_awcache                  : out std_logic_vector(3 downto 0);
    m_axi_wready                   : in  std_logic;
    m_axi_wvalid                   : out std_logic;
    m_axi_wdata                    : out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
    m_axi_wstrb                    : out std_logic_vector((C_M_AXI_DATA_WIDTH)/8 - 1 downto 0);
    m_axi_wlast                    : out std_logic;
    m_axi_bready                   : out std_logic;
    m_axi_bvalid                   : in  std_logic;
    m_axi_bresp                    : in  std_logic_vector(1 downto 0);

    -- Simple Memory Interface:
    mem_go      : in  std_logic;
    mem_clr_go  : out std_logic;
    mem_busy    : out std_logic;
    mem_done    : out std_logic;
    mem_error   : out std_logic;
    mem_timeout : out std_logic;
    
    mem_rd_req      : in std_logic;
    mem_wr_req      : in std_logic;
    mem_bus_lock    : in std_logic;
    mem_burst       : in std_logic;
    mem_addr        : in std_logic_vector(31 downto 0);
    mem_be          : in std_logic_vector(15 downto 0);
    mem_xfer_length : in std_logic_vector(11 downto 0);
    
    mem_in_en   : out std_logic;
    mem_in_data : out std_logic_vector(C_NATIVE_DATA_WIDTH-1 downto 0);

    mem_out_en   : out std_logic;
    mem_out_data : in  std_logic_vector(C_NATIVE_DATA_WIDTH-1 downto 0)
  );

end entity AXI_Master;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture IMP of AXI_Master is

  signal Clk                            : std_logic;
  signal Reset_n                        : std_logic;

  signal mst_cntl_rd_req                : std_logic;
  signal mst_cntl_wr_req                : std_logic;
  signal mst_cntl_bus_lock              : std_logic;
  signal mst_cntl_burst                 : std_logic;
  signal mst_ip2bus_addr                : std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
  signal mst_xfer_length                : std_logic_vector(C_LENGTH_WIDTH-1 downto 0);
  --signal mst_xfer_reg_len               : std_logic_vector(19 downto 0);
  signal mst_ip2bus_be                  : std_logic_vector(15 downto 0);
  signal mst_go                         : std_logic;
  -- signals for master model command interface state machine
  type CMD_CNTL_SM_TYPE is (CMD_IDLE, CMD_RUN, CMD_WAIT_FOR_DATA, CMD_DONE);
  signal mst_cmd_sm_state               : CMD_CNTL_SM_TYPE;
  signal mst_cmd_sm_set_done            : std_logic;
  signal mst_cmd_sm_set_error           : std_logic;
  signal mst_cmd_sm_set_timeout         : std_logic;
  signal mst_cmd_sm_busy                : std_logic;
  signal mst_cmd_sm_clr_go              : std_logic;
  signal mst_cmd_sm_rd_req              : std_logic;
  signal mst_cmd_sm_wr_req              : std_logic;
  signal mst_cmd_sm_reset               : std_logic;
  signal mst_cmd_sm_bus_lock            : std_logic;
  signal mst_cmd_sm_ip2bus_addr         : std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
  signal mst_cmd_sm_ip2bus_be           : std_logic_vector(C_NATIVE_DATA_WIDTH/8-1 downto 0);
  signal mst_cmd_sm_xfer_type           : std_logic;
  signal mst_cmd_sm_xfer_length         : std_logic_vector(C_LENGTH_WIDTH-1 downto 0);
  signal mst_cmd_sm_start_rd_llink      : std_logic;
  signal mst_cmd_sm_start_wr_llink      : std_logic;
  -- signals for master model read locallink interface state machine
  type RD_LLINK_SM_TYPE is (LLRD_IDLE, LLRD_GO);
  signal mst_llrd_sm_state              : RD_LLINK_SM_TYPE;
  signal mst_llrd_sm_dst_rdy            : std_logic;
  -- signals for master model write locallink interface state machine
  type WR_LLINK_SM_TYPE is (LLWR_IDLE, LLWR_SNGL_INIT, LLWR_SNGL, LLWR_BRST_INIT, LLWR_BRST, LLWR_BRST_LAST_BEAT);
  signal mst_llwr_sm_state              : WR_LLINK_SM_TYPE;
  signal mst_llwr_sm_src_rdy            : std_logic;
  signal mst_llwr_sm_sof                : std_logic;
  signal mst_llwr_sm_eof                : std_logic;
  signal mst_llwr_byte_cnt              : integer;
  signal mst_valid_write_xfer           : std_logic;
  signal mst_valid_read_xfer            : std_logic;
  
  -- signals to/from master ipif
  signal ip2bus_mstrd_req               : std_logic;
  signal ip2bus_mstwr_req               : std_logic;
  signal ip2bus_mst_addr                : std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
  signal ip2bus_mst_be                  : std_logic_vector((C_NATIVE_DATA_WIDTH/8)-1 downto 0);
  signal ip2bus_mst_length              : std_logic_vector(C_LENGTH_WIDTH-1 downto 0);
  signal ip2bus_mst_type                : std_logic;
  signal ip2bus_mst_lock                : std_logic;
  signal ip2bus_mst_reset               : std_logic;
  signal bus2ip_mst_cmdack              : std_logic;
  signal bus2ip_mst_cmplt               : std_logic;
  signal bus2ip_mst_error               : std_logic;
  signal bus2ip_mst_rearbitrate         : std_logic;
  signal bus2ip_mst_cmd_timeout         : std_logic;
  signal bus2ip_mstrd_d                 : std_logic_vector(C_NATIVE_DATA_WIDTH-1 downto 0);
  signal bus2ip_mstrd_rem               : std_logic_vector((C_NATIVE_DATA_WIDTH)/8-1 downto 0);
  signal bus2ip_mstrd_sof_n             : std_logic;
  signal bus2ip_mstrd_eof_n             : std_logic;
  signal bus2ip_mstrd_src_rdy_n         : std_logic;
  signal bus2ip_mstrd_src_dsc_n         : std_logic;
  signal ip2bus_mstrd_dst_rdy_n         : std_logic;
  signal ip2bus_mstrd_dst_dsc_n         : std_logic;
  signal ip2bus_mstwr_d                 : std_logic_vector(C_NATIVE_DATA_WIDTH-1 downto 0);
  signal ip2bus_mstwr_rem               : std_logic_vector((C_NATIVE_DATA_WIDTH)/8-1 downto 0);
  signal ip2bus_mstwr_src_rdy_n         : std_logic;
  signal ip2bus_mstwr_src_dsc_n         : std_logic;
  signal ip2bus_mstwr_sof_n             : std_logic;
  signal ip2bus_mstwr_eof_n             : std_logic;
  signal bus2ip_mstwr_dst_rdy_n         : std_logic;
  signal bus2ip_mstwr_dst_dsc_n         : std_logic;
  
  attribute MAX_FANOUT : string;
  attribute SIGIS : string;

  attribute SIGIS of Clk : signal is "CLK";
  attribute SIGIS of Reset_n : signal is "RST";
  attribute SIGIS of ip2bus_mst_reset: signal is "RST";
  
  
  
begin




  ------------------------------------------
  -- Instantiate axi_master_burst
  ------------------------------------------
  AXI_MASTER_BURST_I : entity axi_master_burst_v2_0_7.axi_master_burst
    generic map
    (
      C_M_AXI_ADDR_WIDTH             => C_M_AXI_ADDR_WIDTH,
      C_M_AXI_DATA_WIDTH             => C_M_AXI_DATA_WIDTH,
      C_MAX_BURST_LEN                => C_MAX_BURST_LEN,
      C_NATIVE_DATA_WIDTH            => C_NATIVE_DATA_WIDTH,
      C_LENGTH_WIDTH                 => C_LENGTH_WIDTH,
      C_ADDR_PIPE_DEPTH              => C_ADDR_PIPE_DEPTH,
      C_FAMILY                       => C_FAMILY
    )
    port map
    (
      m_axi_aclk                     => m_axi_aclk,
      m_axi_aresetn                  => m_axi_aresetn,
      md_error                       => md_error,
      m_axi_arready                  => m_axi_arready,
      m_axi_arvalid                  => m_axi_arvalid,
      m_axi_araddr                   => m_axi_araddr,
      m_axi_arlen                    => m_axi_arlen,
      m_axi_arsize                   => m_axi_arsize,
      m_axi_arburst                  => m_axi_arburst,
      m_axi_arprot                   => m_axi_arprot,
      m_axi_arcache                  => m_axi_arcache,
      m_axi_rready                   => m_axi_rready,
      m_axi_rvalid                   => m_axi_rvalid,
      m_axi_rdata                    => m_axi_rdata,
      m_axi_rresp                    => m_axi_rresp,
      m_axi_rlast                    => m_axi_rlast,
      m_axi_awready                  => m_axi_awready,
      m_axi_awvalid                  => m_axi_awvalid,
      m_axi_awaddr                   => m_axi_awaddr,
      m_axi_awlen                    => m_axi_awlen,
      m_axi_awsize                   => m_axi_awsize,
      m_axi_awburst                  => m_axi_awburst,
      m_axi_awprot                   => m_axi_awprot,
      m_axi_awcache                  => m_axi_awcache,
      m_axi_wready                   => m_axi_wready,
      m_axi_wvalid                   => m_axi_wvalid,
      m_axi_wdata                    => m_axi_wdata,
      m_axi_wstrb                    => m_axi_wstrb,
      m_axi_wlast                    => m_axi_wlast,
      m_axi_bready                   => m_axi_bready,
      m_axi_bvalid                   => m_axi_bvalid,
      m_axi_bresp                    => m_axi_bresp,
      ip2bus_mstrd_req               => ip2bus_mstrd_req,
      ip2bus_mstwr_req               => ip2bus_mstwr_req,
      ip2bus_mst_addr                => ip2bus_mst_addr,
      ip2bus_mst_be                  => ip2bus_mst_be,
      ip2bus_mst_length              => ip2bus_mst_length,
      ip2bus_mst_type                => ip2bus_mst_type,
      ip2bus_mst_lock                => ip2bus_mst_lock,
      ip2bus_mst_reset               => ip2bus_mst_reset,
      bus2ip_mst_cmdack              => bus2ip_mst_cmdack,
      bus2ip_mst_cmplt               => bus2ip_mst_cmplt,
      bus2ip_mst_error               => bus2ip_mst_error,
      bus2ip_mst_rearbitrate         => bus2ip_mst_rearbitrate,
      bus2ip_mst_cmd_timeout         => bus2ip_mst_cmd_timeout,
      bus2ip_mstrd_d                 => bus2ip_mstrd_d,
      bus2ip_mstrd_rem               => bus2ip_mstrd_rem,
      bus2ip_mstrd_sof_n             => bus2ip_mstrd_sof_n,
      bus2ip_mstrd_eof_n             => bus2ip_mstrd_eof_n,
      bus2ip_mstrd_src_rdy_n         => bus2ip_mstrd_src_rdy_n,
      bus2ip_mstrd_src_dsc_n         => bus2ip_mstrd_src_dsc_n,
      ip2bus_mstrd_dst_rdy_n         => ip2bus_mstrd_dst_rdy_n,
      ip2bus_mstrd_dst_dsc_n         => ip2bus_mstrd_dst_dsc_n,
      ip2bus_mstwr_d                 => ip2bus_mstwr_d,
      ip2bus_mstwr_rem               => ip2bus_mstwr_rem,
      ip2bus_mstwr_src_rdy_n         => ip2bus_mstwr_src_rdy_n,
      ip2bus_mstwr_src_dsc_n         => ip2bus_mstwr_src_dsc_n,
      ip2bus_mstwr_sof_n             => ip2bus_mstwr_sof_n,
      ip2bus_mstwr_eof_n             => ip2bus_mstwr_eof_n,
      bus2ip_mstwr_dst_rdy_n         => bus2ip_mstwr_dst_rdy_n,
      bus2ip_mstwr_dst_dsc_n         => bus2ip_mstwr_dst_dsc_n
    );


  Clk <= m_axi_aclk;
  Reset_n <= m_axi_aresetn;


  mst_go <= mem_go;
  mem_clr_go <= mst_cmd_sm_clr_go;
  mem_busy <= mst_cmd_sm_busy;
  mem_done <= mst_cmd_sm_set_done;
  mem_error <= mst_cmd_sm_set_error;
  mem_timeout <= mst_cmd_sm_set_timeout;

  mst_cntl_rd_req <= mem_rd_req;
  mst_cntl_wr_req <= mem_wr_req;
  mst_cntl_bus_lock <= mem_bus_lock;
  mst_cntl_burst <= mem_burst;
  mst_ip2bus_addr <= mem_addr;
  mst_ip2bus_be <= mem_be;
  mst_xfer_length <= mem_xfer_length;

  mem_in_en <= mst_valid_read_xfer;
  mem_in_data <= bus2ip_mstrd_d;

  mem_out_en <= mst_valid_write_xfer;
  ip2bus_mstwr_d <= mem_out_data;


  -- user logic master command interface assignments
  IP2Bus_MstRd_Req  <= mst_cmd_sm_rd_req;
  IP2Bus_MstWr_Req  <= mst_cmd_sm_wr_req;
  IP2Bus_Mst_Addr   <= mst_cmd_sm_ip2bus_addr;
  IP2Bus_Mst_BE     <= mst_cmd_sm_ip2bus_be;
  IP2Bus_Mst_Type   <= mst_cmd_sm_xfer_type;
  IP2Bus_Mst_Length <= mst_cmd_sm_xfer_length;
  IP2Bus_Mst_Lock   <= mst_cmd_sm_bus_lock;
  IP2Bus_Mst_Reset  <= mst_cmd_sm_reset;

  --implement master command interface state machine
  MASTER_CMD_SM_PROC : process( Clk ) is
  begin

    if ( Clk'event and Clk = '1' ) then
      if ( Reset_n = '0' ) then

        -- reset condition
        mst_cmd_sm_state          <= CMD_IDLE;
        mst_cmd_sm_clr_go         <= '0';
        mst_cmd_sm_rd_req         <= '0';
        mst_cmd_sm_wr_req         <= '0';
        mst_cmd_sm_bus_lock       <= '0';
        mst_cmd_sm_reset          <= '0';
        mst_cmd_sm_ip2bus_addr    <= (others => '0');
        mst_cmd_sm_ip2bus_be      <= (others => '0');
        mst_cmd_sm_xfer_type      <= '0';
        mst_cmd_sm_xfer_length    <= (others => '0');
        mst_cmd_sm_set_done       <= '0';
        mst_cmd_sm_set_error      <= '0';
        mst_cmd_sm_set_timeout    <= '0';
        mst_cmd_sm_busy           <= '0';
        mst_cmd_sm_start_rd_llink <= '0';
        mst_cmd_sm_start_wr_llink <= '0';


      else

        -- default condition
        mst_cmd_sm_clr_go         <= '0';
        mst_cmd_sm_rd_req         <= '0';
        mst_cmd_sm_wr_req         <= '0';
        mst_cmd_sm_bus_lock       <= '0';
        mst_cmd_sm_reset          <= '0';
        mst_cmd_sm_ip2bus_addr    <= (others => '0');
        mst_cmd_sm_ip2bus_be      <= (others => '0');
        mst_cmd_sm_xfer_type      <= '0';
        mst_cmd_sm_xfer_length    <= (others => '0');
        mst_cmd_sm_set_done       <= '0';
        mst_cmd_sm_set_error      <= '0';
        mst_cmd_sm_set_timeout    <= '0';
        mst_cmd_sm_busy           <= '1';
        mst_cmd_sm_start_rd_llink <= '0';
        mst_cmd_sm_start_wr_llink <= '0';

        -- state transition
        case mst_cmd_sm_state is

          when CMD_IDLE =>
            if ( mst_go = '1' ) then
              mst_cmd_sm_state  <= CMD_RUN;
              mst_cmd_sm_clr_go <= '1';
              if ( mst_cntl_rd_req = '1' ) then
                mst_cmd_sm_start_rd_llink <= '1';
              elsif ( mst_cntl_wr_req = '1' ) then
                mst_cmd_sm_start_wr_llink <= '1';
              end if;
            else
              mst_cmd_sm_state  <= CMD_IDLE;
              mst_cmd_sm_busy   <= '0';
            end if;
            

          when CMD_RUN =>
            if ( Bus2IP_Mst_CmdAck = '1' and Bus2IP_Mst_Cmplt = '0' ) then
              mst_cmd_sm_state <= CMD_WAIT_FOR_DATA;
            elsif ( Bus2IP_Mst_Cmplt = '1' ) then
              mst_cmd_sm_state <= CMD_DONE;
              if ( Bus2IP_Mst_Cmd_Timeout = '1' ) then
                -- AXI4LITE address phase timeout
                mst_cmd_sm_set_error   <= '1';
                mst_cmd_sm_set_timeout <= '1';
              elsif ( Bus2IP_Mst_Error = '1' ) then
                -- AXI4LITE data transfer error
                mst_cmd_sm_set_error   <= '1';
              end if;
            else
              mst_cmd_sm_state       <= CMD_RUN;
              mst_cmd_sm_rd_req      <= mst_cntl_rd_req;
              mst_cmd_sm_wr_req      <= mst_cntl_wr_req;
              mst_cmd_sm_ip2bus_addr <= mst_ip2bus_addr;
              mst_cmd_sm_ip2bus_be   <= mst_ip2bus_be(15 downto 16-C_NATIVE_DATA_WIDTH/8 );
              mst_cmd_sm_xfer_type   <= mst_cntl_burst;
              mst_cmd_sm_xfer_length <= mst_xfer_length;
              mst_cmd_sm_bus_lock    <= mst_cntl_bus_lock;
            end if;
            

          when CMD_WAIT_FOR_DATA =>
            if ( Bus2IP_Mst_Cmplt = '1' ) then
              mst_cmd_sm_state <= CMD_DONE;
              if ( Bus2IP_Mst_Cmd_Timeout = '1' ) then
                -- AXI4LITE address phase timeout
                mst_cmd_sm_set_error   <= '1';
                mst_cmd_sm_set_timeout <= '1';
              elsif ( Bus2IP_Mst_Error = '1' ) then
                -- AXI4LITE data transfer error
                mst_cmd_sm_set_error   <= '1';
              end if;
            else
              mst_cmd_sm_state <= CMD_WAIT_FOR_DATA;
            end if;
            

          when CMD_DONE =>
            mst_cmd_sm_state    <= CMD_IDLE;
            mst_cmd_sm_set_done <= '1';
            mst_cmd_sm_busy     <= '0';
            

          when others =>
            mst_cmd_sm_state    <= CMD_IDLE;
            mst_cmd_sm_busy     <= '0';
            

        end case;

      end if;
    end if;

  end process MASTER_CMD_SM_PROC;

  -- user logic master read locallink interface assignments
  IP2Bus_MstRd_dst_rdy_n <= not(mst_llrd_sm_dst_rdy);
  IP2Bus_MstRd_dst_dsc_n <= '1'; -- do not throttle data

  -- implement a simple state machine to enable the
  -- read locallink interface to transfer data
  LLINK_RD_SM_PROCESS : process( Clk ) is
  begin

    if ( Clk'event and Clk = '1' ) then
      if ( Reset_n = '0' ) then

        -- reset condition
        mst_llrd_sm_state   <= LLRD_IDLE;
        mst_llrd_sm_dst_rdy <= '0';
      else

        -- default condition
        mst_llrd_sm_state   <= LLRD_IDLE;
        mst_llrd_sm_dst_rdy <= '0';

        -- state transition
        case mst_llrd_sm_state is

          when LLRD_IDLE =>
            if ( mst_cmd_sm_start_rd_llink = '1') then
              mst_llrd_sm_state <= LLRD_GO;
            else
              mst_llrd_sm_state <= LLRD_IDLE;
            end if;

          when LLRD_GO =>
            -- done, end of packet
            if ( mst_llrd_sm_dst_rdy    = '1' and
                 Bus2IP_MstRd_src_rdy_n = '0' and
                 Bus2IP_MstRd_eof_n     = '0' ) then
              mst_llrd_sm_state   <= LLRD_IDLE;
            -- not done yet, continue receiving data
            else
              mst_llrd_sm_state   <= LLRD_GO;
              mst_llrd_sm_dst_rdy <= '1';
            end if;

          when others =>
            mst_llrd_sm_state <= LLRD_IDLE;

        end case;

      end if;
    else
      null;
    end if;

  end process LLINK_RD_SM_PROCESS;

  -- user logic master write locallink interface assignments
  IP2Bus_MstWr_src_rdy_n <= not(mst_llwr_sm_src_rdy);
  IP2Bus_MstWr_src_dsc_n <= '1'; -- do not throttle data
  IP2Bus_MstWr_rem       <= (others => '0');
  IP2Bus_MstWr_sof_n     <= not(mst_llwr_sm_sof);
  IP2Bus_MstWr_eof_n     <= not(mst_llwr_sm_eof);

  -- implement a simple state machine to enable the
  -- write locallink interface to transfer data
  LLINK_WR_SM_PROC : process( Clk ) is
    constant BYTES_PER_BEAT : integer := C_NATIVE_DATA_WIDTH/8;
  begin

    if ( Clk'event and Clk = '1' ) then
      if ( Reset_n = '0' ) then

        -- reset condition
        mst_llwr_sm_state   <= LLWR_IDLE;
        mst_llwr_sm_src_rdy <= '0';
        mst_llwr_sm_sof     <= '0';
        mst_llwr_sm_eof     <= '0';
        mst_llwr_byte_cnt   <= 0;
        

      else

        -- default condition
        mst_llwr_sm_state   <= LLWR_IDLE;
        mst_llwr_sm_src_rdy <= '0';
        mst_llwr_sm_sof     <= '0';
        mst_llwr_sm_eof     <= '0';
        mst_llwr_byte_cnt   <= 0;

        -- state transition
        case mst_llwr_sm_state is

          when LLWR_IDLE =>
            if ( mst_cmd_sm_start_wr_llink = '1' and mst_cntl_burst = '0' ) then
              mst_llwr_sm_state <= LLWR_SNGL_INIT;
            elsif ( mst_cmd_sm_start_wr_llink = '1' and mst_cntl_burst = '1' ) then
              mst_llwr_sm_state <= LLWR_BRST_INIT;
            else
              mst_llwr_sm_state <= LLWR_IDLE;
            end if;
            

          when LLWR_SNGL_INIT =>
            mst_llwr_sm_state   <= LLWR_SNGL;
            mst_llwr_sm_src_rdy <= '1';
            mst_llwr_sm_sof     <= '1';
            mst_llwr_sm_eof     <= '1';
            

          when LLWR_SNGL =>
            -- destination discontinue write
            if ( Bus2IP_MstWr_dst_dsc_n = '0' and Bus2IP_MstWr_dst_rdy_n = '0' ) then
              mst_llwr_sm_state   <= LLWR_IDLE;
              mst_llwr_sm_src_rdy <= '0';
              mst_llwr_sm_eof     <= '0';
            -- single data beat transfer complete
            elsif ( mst_valid_write_xfer = '1' ) then
              mst_llwr_sm_state   <= LLWR_IDLE;
              mst_llwr_sm_src_rdy <= '0';
              mst_llwr_sm_sof     <= '0';
              mst_llwr_sm_eof     <= '0';
            -- wait on destination
            else
              mst_llwr_sm_state   <= LLWR_SNGL;
              mst_llwr_sm_src_rdy <= '1';
              mst_llwr_sm_sof     <= '1';
              mst_llwr_sm_eof     <= '1';
            end if;
            

          when LLWR_BRST_INIT =>
            mst_llwr_sm_state   <= LLWR_BRST;
            mst_llwr_sm_src_rdy <= '1';
            mst_llwr_sm_sof     <= '1';
            mst_llwr_byte_cnt   <= CONV_INTEGER(mst_xfer_length);
            
          when LLWR_BRST =>
            if ( mst_valid_write_xfer = '1' ) then
              mst_llwr_sm_sof <= '0';
            else
              mst_llwr_sm_sof <= mst_llwr_sm_sof;
            end if;
            -- destination discontinue write
            if ( Bus2IP_MstWr_dst_dsc_n = '0' and
                 Bus2IP_MstWr_dst_rdy_n = '0' ) then
              mst_llwr_sm_state   <= LLWR_IDLE;
              mst_llwr_sm_src_rdy <= '1';
              mst_llwr_sm_eof     <= '1';
            -- last data beat write
            elsif ( mst_valid_write_xfer = '1' and
                   (mst_llwr_byte_cnt-BYTES_PER_BEAT) <= BYTES_PER_BEAT ) then
              mst_llwr_sm_state   <= LLWR_BRST_LAST_BEAT;
              mst_llwr_sm_src_rdy <= '1';
              mst_llwr_sm_eof     <= '1';
            -- wait on destination
            else
              mst_llwr_sm_state   <= LLWR_BRST;
              mst_llwr_sm_src_rdy <= '1';
              -- decrement write transfer counter if it's a valid write
              if ( mst_valid_write_xfer = '1' ) then
                mst_llwr_byte_cnt <= mst_llwr_byte_cnt - BYTES_PER_BEAT;
              else
                mst_llwr_byte_cnt <= mst_llwr_byte_cnt;
              end if;
            end if;
            

          when LLWR_BRST_LAST_BEAT =>
            -- destination discontinue write
            if ( Bus2IP_MstWr_dst_dsc_n = '0' and
                 Bus2IP_MstWr_dst_rdy_n = '0' ) then
              mst_llwr_sm_state   <= LLWR_IDLE;
              mst_llwr_sm_src_rdy <= '0';
            -- last data beat done
            elsif ( mst_valid_write_xfer = '1' ) then
              mst_llwr_sm_state   <= LLWR_IDLE;
              mst_llwr_sm_src_rdy <= '0';
            -- wait on destination
            else
              mst_llwr_sm_state   <= LLWR_BRST_LAST_BEAT;
              mst_llwr_sm_src_rdy <= '1';
              mst_llwr_sm_eof     <= '1';
            end if;
            

          when others =>
            mst_llwr_sm_state <= LLWR_IDLE;
            

        end case;

      end if;
    else
      null;
    end if;

  end process LLINK_WR_SM_PROC;

  -- local signals 
  mst_valid_read_xfer  <= not(Bus2IP_MstRd_src_rdy_n) and mst_llrd_sm_dst_rdy;
  mst_valid_write_xfer <= not(Bus2IP_MstWr_dst_rdy_n) and mst_llwr_sm_src_rdy;

end IMP;

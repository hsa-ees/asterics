----------------------------------------------------------------------------------
--  This file is part of the ASTERICS Framework.                                  
--  (C) 2019 Hochschule Augsburg, University of Applied Sciences             
----------------------------------------------------------------------------------
-- Entity:         as_canny_pipeline                                                  
--                                                                                
-- Company:        Efficient Embedded Systems Group at                            
--                 University of Applied Sciences, Augsburg, Germany              
-- Author:         as_automatics (automated processing chain generator)           
--                                                                                
-- Modified:                                                                      
--                                                                                
-- Description: ASTERICS module group 'as_canny_pipeline' file generated by Automatics
----------------------------------------------------------------------------------
--  This program is free software; you can redistribute it and/or                 
--  modify it under the terms of the GNU Lesser General Public                    
--  License as published by the Free Software Foundation; either                  
--  version 3 of the License, or (at your option) any later version.              
--                                                                                
--  This program is distributed in the hope that it will be useful,               
--  but WITHOUT ANY WARRANTY; without even the implied warranty of                
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU             
--  Lesser General Public License for more details.                               
--                                                                                
--  You should have received a copy of the GNU Lesser General Public License      
--  along with this program; if not, see <http://www.gnu.org/licenses/>           
--  or write to the Free Software Foundation, Inc.,                               
--  51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.                 
----------------------------------------------------------------------------------
--! @file  as_canny_pipeline.vhd
--! @brief Canny edge detector implementation generated using Automatics.
--! @addtogroup asterics_modules
--! @{
--! @defgroup as_canny_pipeline as_canny_pipeline: Canny Edge Detector
--! Canny edge detector implementation using ASTERICS modules and the
--! 2D Window Pipeline architecture.
--! Original design by Markus Bihler, Automatics compatible design by Philip Manke.
--! @}
----------------------------------------------------------------------------------

--! @addtogroup as_canny_pipeline
--! @{

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library asterics;
use asterics.helpers.all;
use asterics.as_generic_filter.all;
use asterics.as_2d_conv_filter_internal;
use asterics.as_cordic_direction;
use asterics.as_edge_list;
use asterics.as_edge_nms;
use asterics.as_edge_threshold;
use asterics.as_feature_counter;
use asterics.as_gradient_weight;
use asterics.as_pipeline_flush;
use asterics.as_pipeline_row;

entity as_canny_pipeline is
  generic(
    DIN_WIDTH : integer := 8;
    LINE_WIDTH : integer := 640;
    IMAGE_HEIGHT : integer := 480;
    MINIMUM_BRAM_SIZE : integer := 256
  );
  port(
    reset : in std_logic;
    clk : in std_logic;
    slv_reg_config : out slv_reg_config_table(0 to 4);
    slv_ctrl_reg : in slv_reg_data(0 to 4);
    slv_status_reg : out slv_reg_data(0 to 4);
    slv_reg_modify : out std_logic_vector(0 to 4);
    cam0_vsync : in std_logic;
    cam0_hsync : in std_logic;
    cam0_strobe : in std_logic;
    cam0_data : in std_logic_vector(7 downto 0);
    cam0_vcomplete : in std_logic;
    cam0_data_error : in std_logic;
    cam0_stall : out std_logic;
    feat_strobe : out std_logic;
    feat_data : out std_logic_vector(31 downto 0);
    feat_data_unit_complete : out std_logic
  );
end entity as_canny_pipeline;

--! @}

architecture RTL of as_canny_pipeline is

  -- Constant declarations:
  constant slave_register_configuration : slv_reg_config_table(0 to 4) := (AS_REG_BOTH, AS_REG_STATUS, AS_REG_CONTROL, AS_REG_NONE, AS_REG_STATUS);
  -- Glue signals:
  signal fsobelx_data_out : std_logic_vector(8 downto 0);
  signal fsobely_data_out : std_logic_vector(8 downto 0);
  signal cordic_data_out_reduced : std_logic_vector(1 downto 0);
  signal nms_data_out : std_logic_vector(8 downto 0);
  signal thresh_data_out : std_logic_vector(1 downto 0);
  signal cordic_data_out_full : std_logic_vector(10 downto 0);
  signal reset_int : std_logic;
  signal flush_done_int : std_logic;
  signal flush : std_logic;
  signal ready : std_logic;
  signal strobe_int_out : std_logic;
  signal strobe_int : std_logic;
  signal stall_out_int : std_logic;
  signal sw_reset : std_logic;
  signal data_stream_in : std_logic_vector(9 downto 0);
  signal pipeline_stream_in : std_logic_vector(9 downto 0);
  signal result_stream_out : std_logic_vector(31 downto 0);
  signal data_stream_out : std_logic_vector(31 downto 0);
  signal reg_modify_vect : std_logic_vector(0 to 4);
  signal s_register_id0 : std_logic_vector(31 downto 0);
  signal s_register_id1 : std_logic_vector(31 downto 0);
  signal thr_low_in_signal : std_logic_vector(7 downto 0);
  signal s_register_id2 : std_logic_vector(31 downto 0);
  signal thr_high_in_signal : std_logic_vector(7 downto 0);
  signal s_register_id4 : std_logic_vector(31 downto 0);
  signal cam0_data_stream_in : std_logic_vector(7 downto 0);
  signal cam0_hsync_stream_in : std_logic;
  signal cam0_vsync_stream_in : std_logic;
  signal feat_data_out_synced : std_logic_vector(31 downto 0);
  signal cordic_data_out_reduced_delay_input_0 : std_logic_vector(1 downto 0);
  signal cordic_data_out_reduced_delayed_0 : std_logic_vector(1 downto 0);
  signal cordic_data_out_full_delay_input_0 : std_logic_vector(10 downto 0);
  signal cordic_data_out_full_delayed_0 : std_logic_vector(10 downto 0);
  signal cam0_vsync_stream_in_delay_input_0 : std_logic;
  signal cam0_vsync_stream_in_delayed_0 : std_logic;
  signal cam0_hsync_stream_in_delay_input_0 : std_logic;
  signal cam0_hsync_stream_in_delayed_0 : std_logic;
  signal fgauss0_row_0 : std_logic_vector(7 downto 0);
  signal fgauss0_row_1 : std_logic_vector(7 downto 0);
  signal fgauss0_row_2 : std_logic_vector(7 downto 0);
  signal fgauss0_row_3 : std_logic_vector(7 downto 0);
  signal fgauss0_row_4 : std_logic_vector(7 downto 0);
  signal fsobelx_row_0 : std_logic_vector(7 downto 0);
  signal fsobelx_row_1 : std_logic_vector(7 downto 0);
  signal fsobelx_row_2 : std_logic_vector(7 downto 0);
  signal nms_row_0 : std_logic_vector(8 downto 0);
  signal nms_row_1 : std_logic_vector(8 downto 0);
  signal nms_row_2 : std_logic_vector(8 downto 0);
  signal thresh_row_0 : std_logic_vector(1 downto 0);
  signal thresh_row_1 : std_logic_vector(1 downto 0);
  signal strobe_in_combined : std_logic;
  signal feat_data_out_signal : std_logic_vector(31 downto 0);
  signal strobe_out_fixed_value : std_logic;
  signal stall_in_combined : std_logic;
  signal cordic_data_out_full_delay_input_0_intermediate : std_logic_vector(10 downto 0);
  signal cam0_vsync_stream_in_delayed_loopdelay_0 : std_logic;
  signal cam0_vsync_stream_in_delayed_0_last_delay : std_logic;
  signal cam0_hsync_stream_in_delayed_loopdelay_0 : std_logic;
  signal cam0_hsync_stream_in_delayed_0_last_delay : std_logic;
  signal cordic_out_reduced_buffer_line_0_data_in : std_logic_vector(12 downto 0);
  signal cordic_reduced_buffer_line_0_data_out : std_logic_vector(12 downto 0);
  signal cordic_out_reduced_buffer_0_line_data : t_generic_line(0 to 0, 12 downto 0);
  signal cordic_out_full_buffer_line_0_data_in : std_logic_vector(10 downto 0);
  signal cordic_full_buffer_line_0_data_out : std_logic_vector(10 downto 0);
  signal cordic_out_full_buffer_0_line_data : t_generic_line(0 to 0, 10 downto 0);
  signal as_canny_pipeline_cam0_vsync_stream_buffer_line_0_data_in : std_logic_vector(3 downto 0);
  signal as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_data_out : std_logic_vector(3 downto 0);
  signal as_canny_pipeline_cam0_vsync_stream_in_buffer_0_line_data : t_generic_line(0 to 0, 3 downto 0);
  signal cam0_stream_buffer_row_0_data_in : std_logic_vector(67 downto 0);
  signal cam0_stream_in_buffer_row_0_data_out : std_logic_vector(67 downto 0);
  signal fgauss0_data_out_signal : std_logic_vector(7 downto 0);
  signal edge_weight_data_out_signal : std_logic_vector(8 downto 0);
  signal cam0_stream_in_buffer_row_0_line_data : t_generic_line(0 to 4, 67 downto 0);
  signal cam0_stream_buffer_row_4_end_data_in : std_logic_vector(7 downto 0);
  signal cam0_stream_in_buffer_row_4_end_data_out : std_logic_vector(7 downto 0);
  signal cam0_stream_in_buffer_row_4_end_line_data : t_generic_line(0 to 4, 7 downto 0);
  signal fgauss0_buffer_row_2_end_data_in : std_logic_vector(18 downto 0);
  signal fgauss0_buffer_row_2_end_data_out : std_logic_vector(18 downto 0);
  signal fgauss0_buffer_row_2_end_line_data : t_generic_line(0 to 2, 18 downto 0);
  signal as_canny_pipeline_cam0_vsync_stream_buffer_line_0_last_delay_data_in : std_logic_vector(1 downto 0);
  signal as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_last_delay_data_out : std_logic_vector(1 downto 0);
  signal as_canny_pipeline_cam0_vsync_stream_in_buffer_0_last_delay_line_data : t_generic_line(0 to 0, 1 downto 0);
  signal fgauss0_window_in : t_generic_window(0 to 4, 0 to 4, 7 downto 0);
  signal fsobelx_window_in : t_generic_window(0 to 2, 0 to 2, 7 downto 0);
  signal fsobely_window_in : t_generic_window(0 to 2, 0 to 2, 7 downto 0);
  signal nms_window_in : t_generic_window(0 to 2, 0 to 2, 8 downto 0);
  signal thresh_window_in : t_generic_window(0 to 2, 0 to 1, 1 downto 0);
  signal feat_strobe_out_signal : std_logic;
begin

  -- Register assignments:
  slv_reg_config <= slave_register_configuration;
  slv_reg_modify <= reg_modify_vect;
  s_register_id0 <= slv_ctrl_reg(0);
  s_register_id2 <= slv_ctrl_reg(2);
  slv_status_reg(1) <= s_register_id1;
  slv_status_reg(4) <= s_register_id4;

  -- Assigning window signals:
  assign_windows_p : process(strobe_int, cam0_stream_in_buffer_row_0_line_data, cam0_stream_in_buffer_row_4_end_line_data, fgauss0_buffer_row_2_end_line_data) is
  begin
    -- Build window 'fgauss0_window_in'
    f_set_line_of_generic_window(fgauss0_window_in, 0, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 0, 8));
    f_set_line_of_generic_window(fgauss0_window_in, 1, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 8, 8));
    f_set_line_of_generic_window(fgauss0_window_in, 2, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 16, 8));
    f_set_line_of_generic_window(fgauss0_window_in, 3, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 24, 8));
    f_set_line_of_generic_window(fgauss0_window_in, 4, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_4_end_line_data, 0, 8));
  
    -- Build window 'fsobelx_window_in'
    f_set_line_of_generic_window(fsobelx_window_in, 0, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 32, 8));
    f_set_line_of_generic_window(fsobelx_window_in, 1, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 40, 8));
    f_set_line_of_generic_window(fsobelx_window_in, 2, f_cut_vectors_of_generic_line(fgauss0_buffer_row_2_end_line_data, 0, 8));
  
    -- Build window 'fsobely_window_in'
    f_set_line_of_generic_window(fsobely_window_in, 0, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 32, 8));
    f_set_line_of_generic_window(fsobely_window_in, 1, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 40, 8));
    f_set_line_of_generic_window(fsobely_window_in, 2, f_cut_vectors_of_generic_line(fgauss0_buffer_row_2_end_line_data, 0, 8));
  
    -- Build window 'nms_window_in'
    f_set_line_of_generic_window(nms_window_in, 0, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 48, 9));
    f_set_line_of_generic_window(nms_window_in, 1, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 57, 9));
    f_set_line_of_generic_window(nms_window_in, 2, f_cut_vectors_of_generic_line(fgauss0_buffer_row_2_end_line_data, 8, 9));
  
    -- Build window 'thresh_window_in'
    f_set_line_of_generic_window(thresh_window_in, 0, f_cut_vectors_of_generic_line(cam0_stream_in_buffer_row_0_line_data, 66, 2));
    f_set_line_of_generic_window(thresh_window_in, 1, f_cut_vectors_of_generic_line(fgauss0_buffer_row_2_end_line_data, 17, 2));
  
  end process;

  
  -- Port assignments:
  

  -- Bundled signals:
  
  -- Signal assignments:
  reset_int <= reset or sw_reset;
  feat_data_unit_complete <= flush_done_int;
  cam0_stall <= stall_out_int;

  -- Assign to signal data_stream_in:
  data_stream_in(7 downto 0) <= cam0_data;
  data_stream_in(8) <= cam0_hsync;
  data_stream_in(9) <= cam0_vsync;


  -- Assign from signal pipeline_stream_in:
  cam0_data_stream_in <= pipeline_stream_in(7 downto 0);
  cam0_hsync_stream_in <= pipeline_stream_in(8);
  cam0_vsync_stream_in <= pipeline_stream_in(9);


  -- Assign to signal result_stream_out:
  result_stream_out(31 downto 0) <= feat_data_out_signal;


  -- Assign from signal data_stream_out:
  feat_data_out_synced <= data_stream_out(31 downto 0);


  -- Assign to signal reg_modify_vect:
  reg_modify_vect(0) <= '-';
  reg_modify_vect(1) <= '1';
  reg_modify_vect(2) <= '0';
  reg_modify_vect(3) <= '0';
  reg_modify_vect(4) <= '1';


  -- Assign from signal s_register_id0:
  sw_reset <= s_register_id0(0);
  flush <= s_register_id0(1);


  -- Assign to signal s_register_id1:
  s_register_id1(0) <= ready;
  s_register_id1(31 downto 1) <= (others => '0');


  -- Assign from signal s_register_id2:
  thr_low_in_signal <= s_register_id2(7 downto 0);
  thr_high_in_signal <= s_register_id2(15 downto 8);

  cam0_hsync_stream_in_delay_input_0 <= cam0_hsync_stream_in;
  cam0_vsync_stream_in_delay_input_0 <= cam0_vsync_stream_in;
  feat_data <= feat_data_out_synced;
  strobe_in_combined <= cam0_strobe;
  feat_strobe <= strobe_out_fixed_value;
  strobe_out_fixed_value <= strobe_int_out and feat_strobe_out_signal;

  -- Assign to signal cordic_out_reduced_buffer_line_0_data_in:
  cordic_out_reduced_buffer_line_0_data_in(1 downto 0) <= cordic_data_out_reduced_delay_input_0;
  cordic_out_reduced_buffer_line_0_data_in(12 downto 2) <= cordic_data_out_full_delay_input_0;


  -- Assign from signal cordic_reduced_buffer_line_0_data_out:
  cordic_data_out_reduced_delayed_0 <= cordic_reduced_buffer_line_0_data_out(1 downto 0);
  cordic_data_out_full_delay_input_0_intermediate <= cordic_reduced_buffer_line_0_data_out(12 downto 2);


  -- Assign to signal cordic_out_full_buffer_line_0_data_in:
  cordic_out_full_buffer_line_0_data_in(10 downto 0) <= cordic_data_out_full_delay_input_0_intermediate;


  -- Assign from signal cordic_full_buffer_line_0_data_out:
  cordic_data_out_full_delayed_0 <= cordic_full_buffer_line_0_data_out(10 downto 0);


  -- Assign to signal as_canny_pipeline_cam0_vsync_stream_buffer_line_0_data_in:
  as_canny_pipeline_cam0_vsync_stream_buffer_line_0_data_in(0) <= cam0_vsync_stream_in_delay_input_0;
  as_canny_pipeline_cam0_vsync_stream_buffer_line_0_data_in(1) <= cam0_vsync_stream_in_delayed_loopdelay_0;
  as_canny_pipeline_cam0_vsync_stream_buffer_line_0_data_in(2) <= cam0_hsync_stream_in_delay_input_0;
  as_canny_pipeline_cam0_vsync_stream_buffer_line_0_data_in(3) <= cam0_hsync_stream_in_delayed_loopdelay_0;


  -- Assign from signal as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_data_out:
  cam0_vsync_stream_in_delayed_loopdelay_0 <= as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_data_out(0);
  cam0_vsync_stream_in_delayed_0_last_delay <= as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_data_out(1);
  cam0_hsync_stream_in_delayed_loopdelay_0 <= as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_data_out(2);
  cam0_hsync_stream_in_delayed_0_last_delay <= as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_data_out(3);


  -- Assign to signal cam0_stream_buffer_row_0_data_in:
  cam0_stream_buffer_row_0_data_in(7 downto 0) <= cam0_data_stream_in;
  cam0_stream_buffer_row_0_data_in(15 downto 8) <= fgauss0_row_0;
  cam0_stream_buffer_row_0_data_in(23 downto 16) <= fgauss0_row_1;
  cam0_stream_buffer_row_0_data_in(31 downto 24) <= fgauss0_row_2;
  cam0_stream_buffer_row_0_data_in(39 downto 32) <= fgauss0_data_out_signal;
  cam0_stream_buffer_row_0_data_in(47 downto 40) <= fsobelx_row_0;
  cam0_stream_buffer_row_0_data_in(56 downto 48) <= edge_weight_data_out_signal;
  cam0_stream_buffer_row_0_data_in(65 downto 57) <= nms_row_0;
  cam0_stream_buffer_row_0_data_in(67 downto 66) <= thresh_data_out;


  -- Assign from signal cam0_stream_in_buffer_row_0_data_out:
  fgauss0_row_0 <= cam0_stream_in_buffer_row_0_data_out(7 downto 0);
  fgauss0_row_1 <= cam0_stream_in_buffer_row_0_data_out(15 downto 8);
  fgauss0_row_2 <= cam0_stream_in_buffer_row_0_data_out(23 downto 16);
  fgauss0_row_3 <= cam0_stream_in_buffer_row_0_data_out(31 downto 24);
  fsobelx_row_0 <= cam0_stream_in_buffer_row_0_data_out(39 downto 32);
  fsobelx_row_1 <= cam0_stream_in_buffer_row_0_data_out(47 downto 40);
  nms_row_0 <= cam0_stream_in_buffer_row_0_data_out(56 downto 48);
  nms_row_1 <= cam0_stream_in_buffer_row_0_data_out(65 downto 57);
  thresh_row_0 <= cam0_stream_in_buffer_row_0_data_out(67 downto 66);


  -- Assign to signal cam0_stream_buffer_row_4_end_data_in:
  cam0_stream_buffer_row_4_end_data_in(7 downto 0) <= fgauss0_row_3;


  -- Assign from signal cam0_stream_in_buffer_row_4_end_data_out:
  fgauss0_row_4 <= cam0_stream_in_buffer_row_4_end_data_out(7 downto 0);


  -- Assign to signal fgauss0_buffer_row_2_end_data_in:
  fgauss0_buffer_row_2_end_data_in(7 downto 0) <= fsobelx_row_1;
  fgauss0_buffer_row_2_end_data_in(16 downto 8) <= nms_row_1;
  fgauss0_buffer_row_2_end_data_in(18 downto 17) <= thresh_row_0;


  -- Assign from signal fgauss0_buffer_row_2_end_data_out:
  fsobelx_row_2 <= fgauss0_buffer_row_2_end_data_out(7 downto 0);
  nms_row_2 <= fgauss0_buffer_row_2_end_data_out(16 downto 8);
  thresh_row_1 <= fgauss0_buffer_row_2_end_data_out(18 downto 17);


  -- Assign to signal as_canny_pipeline_cam0_vsync_stream_buffer_line_0_last_delay_data_in:
  as_canny_pipeline_cam0_vsync_stream_buffer_line_0_last_delay_data_in(0) <= cam0_vsync_stream_in_delayed_0_last_delay;
  as_canny_pipeline_cam0_vsync_stream_buffer_line_0_last_delay_data_in(1) <= cam0_hsync_stream_in_delayed_0_last_delay;


  -- Assign from signal as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_last_delay_data_out:
  cam0_vsync_stream_in_delayed_0 <= as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_last_delay_data_out(0);
  cam0_hsync_stream_in_delayed_0 <= as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_last_delay_data_out(1);

  
  -- Components:

  -- Instantiate module as_pipeline_flush_0:
  as_pipeline_flush_0 : entity as_pipeline_flush
  generic map(
    DIN_WIDTH => 10,
    DOUT_WIDTH => 32,
    PIPELINE_DEPTH => 2574,
    IS_FLUSHDATA_CONSTANT => True,
    CONSTANT_DATA_VALUE => 128
  )
  port map(
    ready => ready,
    flush_done_out => flush_done_int,
    result_data_in => result_stream_out,
    clk => clk,
    reset => reset_int,
    flush_in => flush,
    input_strobe_in => strobe_in_combined,
    input_data_in => data_stream_in,
    input_stall_out => stall_out_int,
    pipeline_strobe_out => strobe_int,
    pipeline_data_out => pipeline_stream_in,
    output_stall_in => stall_in_combined,
    output_strobe_out => strobe_int_out,
    output_data_out => data_stream_out
  );


  -- Instantiate module fgauss0:
  fgauss0 : entity as_2d_conv_filter_internal
  port map(
    data_out => fgauss0_data_out_signal,
    clk => clk,
    reset => reset_int,
    strobe_in => strobe_int,
    window_in => fgauss0_window_in
  );


  -- Instantiate module fsobelx:
  fsobelx : entity as_2d_conv_filter_internal
  generic map(
    DOUT_WIDTH => 9,
    KERNEL_SIZE => 3,
    KERNEL_TYPE => "sobel_x",
    OUTPUT_SIGNED => true
  )
  port map(
    data_out => fsobelx_data_out,
    clk => clk,
    reset => reset_int,
    strobe_in => strobe_int,
    window_in => fsobelx_window_in
  );


  -- Instantiate module fsobely:
  fsobely : entity as_2d_conv_filter_internal
  generic map(
    DOUT_WIDTH => 9,
    KERNEL_SIZE => 3,
    KERNEL_TYPE => "sobel_y",
    OUTPUT_SIGNED => true
  )
  port map(
    data_out => fsobely_data_out,
    clk => clk,
    reset => reset_int,
    strobe_in => strobe_int,
    window_in => fsobely_window_in
  );


  -- Instantiate module edge_weight:
  edge_weight : entity as_gradient_weight
  generic map(
    DIN_WIDTH => 9
  )
  port map(
    data1_in => fsobelx_data_out,
    data2_in => fsobely_data_out,
    data_out => edge_weight_data_out_signal,
    clk => clk,
    reset => reset_int,
    strobe_in => strobe_int
  );


  -- Instantiate module cordic:
  cordic : entity as_cordic_direction
  generic map(
    DIN_WIDTH => 9,
    CORDIC_STEP_COUNT => 9,
    ANGLE_WIDTH => 10
  )
  port map(
    data_x_in => fsobelx_data_out,
    data_y_in => fsobely_data_out,
    data_out_reduced => cordic_data_out_reduced_delay_input_0,
    data_out_full => cordic_data_out_full_delay_input_0,
    clk => clk,
    reset => reset_int,
    strobe_in => strobe_int
  );


  -- Instantiate module nms:
  nms : entity as_edge_nms
  port map(
    data_dir_in => cordic_data_out_reduced_delayed_0,
    data_out => nms_data_out,
    clk => clk,
    reset => reset_int,
    strobe_in => strobe_int,
    window_weight_in => nms_window_in
  );


  -- Instantiate module thresh:
  thresh : entity as_edge_threshold
  port map(
    nms_in => nms_data_out,
    thr_low_in => thr_low_in_signal,
    thr_high_in => thr_high_in_signal,
    data_out => thresh_data_out,
    clk => clk,
    reset => reset_int,
    strobe_in => strobe_int,
    first_row_is_edge => thresh_window_in
  );


  -- Instantiate module feat:
  feat : entity as_edge_list
  generic map(
    DIN_WIDTH => 11,
    X_COORDINATE_WIDTH => 10,
    Y_COORDINATE_WIDTH => 10
  )
  port map(
    is_edge_in => thresh_data_out,
    vsync_in => cam0_vsync_stream_in_delayed_0,
    hsync_in => cam0_hsync_stream_in_delayed_0,
    edge_data_in => cordic_data_out_full_delayed_0,
    clk => clk,
    reset => reset_int,
    strobe_in => strobe_int,
    strobe_out => feat_strobe_out_signal,
    data_out => feat_data_out_signal
  );


  -- Instantiate module featcount:
  featcount : entity as_feature_counter
  port map(
    trigger_in => strobe_out_fixed_value,
    frame_done => flush_done_int,
    count_out => s_register_id4,
    clk => clk,
    reset => reset_int
  );


  -- Instantiate module cordic_data_out_reduced_buffer_line_0:
  cordic_data_out_reduced_buffer_line_0 : entity as_pipeline_row
  generic map(
    DATA_WIDTH => 13,
    WINDOW_WIDTH => 1,
    LINE_WIDTH => 632,
    MINIMUM_LENGTH_FOR_BRAM => 500
  )
  port map(
    buff_in => cordic_out_reduced_buffer_line_0_data_in,
    line_out => cordic_out_reduced_buffer_0_line_data,
    data_out => cordic_reduced_buffer_line_0_data_out,
    clk => clk,
    reset => reset_int,
    strobe => strobe_int
  );


  -- Instantiate module cordic_data_out_full_buffer_line_0:
  cordic_data_out_full_buffer_line_0 : entity as_pipeline_row
  generic map(
    DATA_WIDTH => 11,
    WINDOW_WIDTH => 1,
    LINE_WIDTH => 2,
    MINIMUM_LENGTH_FOR_BRAM => 500
  )
  port map(
    buff_in => cordic_out_full_buffer_line_0_data_in,
    line_out => cordic_out_full_buffer_0_line_data,
    data_out => cordic_full_buffer_line_0_data_out,
    clk => clk,
    reset => reset_int,
    strobe => strobe_int
  );


  -- Instantiate module as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0:
  as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0 : entity as_pipeline_row
  generic map(
    DATA_WIDTH => 4,
    WINDOW_WIDTH => 1,
    LINE_WIDTH => 1286,
    MINIMUM_LENGTH_FOR_BRAM => 500
  )
  port map(
    buff_in => as_canny_pipeline_cam0_vsync_stream_buffer_line_0_data_in,
    line_out => as_canny_pipeline_cam0_vsync_stream_in_buffer_0_line_data,
    data_out => as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_data_out,
    clk => clk,
    reset => reset_int,
    strobe => strobe_int
  );


  -- Instantiate module cam0_data_stream_in_buffer_row_0:
  cam0_data_stream_in_buffer_row_0 : entity as_pipeline_row
  generic map(
    DATA_WIDTH => 68,
    WINDOW_WIDTH => 5,
    LINE_WIDTH => 640,
    MINIMUM_LENGTH_FOR_BRAM => 500
  )
  port map(
    buff_in => cam0_stream_buffer_row_0_data_in,
    line_out => cam0_stream_in_buffer_row_0_line_data,
    data_out => cam0_stream_in_buffer_row_0_data_out,
    clk => clk,
    reset => reset_int,
    strobe => strobe_int
  );


  -- Instantiate module cam0_data_stream_in_buffer_row_4_end:
  cam0_data_stream_in_buffer_row_4_end : entity as_pipeline_row
  generic map(
    DATA_WIDTH => 8,
    WINDOW_WIDTH => 5,
    LINE_WIDTH => 5,
    MINIMUM_LENGTH_FOR_BRAM => 500
  )
  port map(
    buff_in => cam0_stream_buffer_row_4_end_data_in,
    line_out => cam0_stream_in_buffer_row_4_end_line_data,
    data_out => cam0_stream_in_buffer_row_4_end_data_out,
    clk => clk,
    reset => reset_int,
    strobe => strobe_int
  );


  -- Instantiate module fgauss0_buffer_row_2_end:
  fgauss0_buffer_row_2_end : entity as_pipeline_row
  generic map(
    DATA_WIDTH => 19,
    WINDOW_WIDTH => 3,
    LINE_WIDTH => 3,
    MINIMUM_LENGTH_FOR_BRAM => 500
  )
  port map(
    buff_in => fgauss0_buffer_row_2_end_data_in,
    line_out => fgauss0_buffer_row_2_end_line_data,
    data_out => fgauss0_buffer_row_2_end_data_out,
    clk => clk,
    reset => reset_int,
    strobe => strobe_int
  );


  -- Instantiate module as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_last_delay:
  as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_last_delay : entity as_pipeline_row
  generic map(
    DATA_WIDTH => 2,
    WINDOW_WIDTH => 1,
    LINE_WIDTH => 1,
    MINIMUM_LENGTH_FOR_BRAM => 500
  )
  port map(
    buff_in => as_canny_pipeline_cam0_vsync_stream_buffer_line_0_last_delay_data_in,
    line_out => as_canny_pipeline_cam0_vsync_stream_in_buffer_0_last_delay_line_data,
    data_out => as_canny_pipeline_cam0_vsync_stream_in_buffer_line_0_last_delay_data_out,
    clk => clk,
    reset => reset_int,
    strobe => strobe_int
  );

end architecture RTL;
